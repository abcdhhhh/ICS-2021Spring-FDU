`ifndef __MYCPU_DEFS_SVH__
`define __MYCPU_DEFS_SVH__

`include "common.svh"

`include "instr.svh"
`include "cp0.svh"
`include "type.svh"

`endif
